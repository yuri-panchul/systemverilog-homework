`define PD(SYMBOL) $sformatf("SYMBOL:%d", SYMBOL)
`define PB(SYMBOL) $sformatf("SYMBOL:%b", SYMBOL)
`define PH(SYMBOL) $sformatf("SYMBOL:%h", SYMBOL)
